module sieve (clk, rst, in$din, out$wr, out$done, out$addr, out$rdy, out$dout);
    input clk;
    input rst;
    input [7:0] in$din;
    output out$wr;
    output out$done;
    output [7:0] out$addr;
    output out$rdy;
    output [7:0] out$dout;
    reg reg$wr$5;
    reg [7:0] reg$dout$10;
    reg [7:0] reg$addr$15;
    reg reg$rdy$19;
    reg reg$done$23;
    reg [7:0] reg$i$43;
    reg [7:0] reg$end$76;
    assign out$wr = reg$wr$5;
    assign out$done = reg$done$23;
    assign out$addr = reg$addr$15;
    assign out$rdy = reg$rdy$19;
    assign out$dout = reg$dout$10;
    wire [7:0] _$0 = in$din;
    wire _$6 = reg$wr$5;
    wire _$7 = 1'b0;
    wire [7:0] _$11 = reg$dout$10;
    wire [7:0] _$12 = 8'd0;
    wire [7:0] _$16 = reg$addr$15;
    wire _$20 = reg$rdy$19;
    wire _$24 = reg$done$23;
    wire _$28 = 1'b1;
    wire [7:0] _$31 = 8'd100;
    wire _$32 = (_$16 <= _$31);
    wire [7:0] _$40 = 8'd1;
    wire [7:0] _$41 = (_$16 + _$40);
    wire [7:0] _$44 = reg$i$43;
    wire [7:0] _$45 = 8'd2;
    wire _$48 = (_$44 <= _$31);
    wire [7:0] _$52 = (_$44 + _$44);
    wire [7:0] _$64 = (_$16 + _$44);
    wire [7:0] _$73 = (_$44 + _$40);
    wire [7:0] _$77 = reg$end$76;
    wire _$94 = (! _$0);
    wire [7:0] _$104 = (_$77 + _$40);
    wire _$109 = (_$16 < _$77);
    wire _$126 = (_$41 <= _$31);
    wire _$127 = (_$28 && _$126);
    wire _$128 = (! _$126);
    wire _$129 = (_$28 && _$128);
    wire _$130 = (_$28 && _$94);
    wire _$131 = (! _$94);
    wire _$132 = (_$28 && _$131);
    wire _$133 = (_$64 <= _$31);
    wire _$134 = (_$28 && _$133);
    wire _$135 = (! _$133);
    wire _$136 = (_$28 && _$135);
    wire _$137 = (_$73 <= _$31);
    wire _$138 = (_$28 && _$137);
    wire _$139 = (_$132 && _$137);
    wire _$140 = (! _$137);
    wire _$141 = (_$28 && _$140);
    wire _$142 = (_$132 && _$140);
    wire _$143 = (_$136 && _$137);
    wire _$144 = (_$136 && _$140);
    wire [7:0] _$145 = (_$45 + _$45);
    wire [7:0] _$146 = (_$73 + _$73);
    wire _$147 = (_$145 <= _$31);
    wire _$148 = (_$129 && _$147);
    wire _$149 = (_$146 <= _$31);
    wire _$150 = (_$138 && _$149);
    wire _$151 = (_$143 && _$149);
    wire _$152 = (! _$147);
    wire _$153 = (_$129 && _$152);
    wire _$154 = (! _$149);
    wire _$155 = (_$138 && _$154);
    wire _$156 = (_$143 && _$154);
    wire _$157 = (_$41 < _$77);
    wire _$158 = (_$28 && _$157);
    wire _$159 = (_$12 < _$104);
    wire _$160 = (_$141 && _$159);
    wire _$161 = (_$12 < _$77);
    wire _$162 = (_$142 && _$161);
    wire _$163 = (! _$157);
    wire _$164 = (_$28 && _$163);
    wire _$165 = (! _$159);
    wire _$166 = (_$141 && _$165);
    wire _$167 = (! _$161);
    wire _$168 = (_$142 && _$167);
    wire _$169 = (_$151 || _$134);
    wire [7:0] _$170 = (_$151 ? _$146 : _$64);
    wire [7:0] _$171 = (_$151 ? _$73 : _$44);
    wire _$172 = (_$158 || _$164);
    wire [7:0] _$173 = (_$158 ? _$41 : _$41);
    wire _$174 = (_$158 ? _$24 : _$28);
    wire _$175 = (_$160 || _$138);
    wire [7:0] _$176 = (_$160 ? _$12 : _$73);
    wire [7:0] _$177 = (_$160 ? _$73 : _$73);
    wire [7:0] _$178 = (_$160 ? _$104 : _$104);
    wire _$179 = (_$160 ? _$28 : _$20);
    wire _$180 = (_$160 ? _$7 : _$7);
    wire _$181 = (_$175 || _$166);
    wire [7:0] _$182 = (_$175 ? _$176 : _$12);
    wire [7:0] _$183 = (_$175 ? _$177 : _$73);
    wire [7:0] _$184 = (_$175 ? _$178 : _$104);
    wire _$185 = (_$175 ? _$179 : _$28);
    wire _$186 = (_$175 ? _$24 : _$28);
    wire _$187 = (_$175 ? _$180 : _$7);
    wire _$188 = (_$127 || _$153);
    wire [7:0] _$189 = (_$127 ? _$41 : _$145);
    wire [7:0] _$190 = (_$127 ? _$11 : _$40);
    wire [7:0] _$191 = (_$127 ? _$44 : _$45);
    wire _$192 = (_$127 ? _$6 : _$7);
    wire _$193 = (_$188 || _$148);
    wire [7:0] _$194 = (_$188 ? _$189 : _$145);
    wire [7:0] _$195 = (_$188 ? _$190 : _$40);
    wire [7:0] _$196 = (_$188 ? _$191 : _$45);
    wire _$197 = (_$188 ? _$192 : _$6);
    wire _$198 = (_$155 || _$141);
    wire [7:0] _$199 = (_$155 ? _$146 : _$45);
    wire [7:0] _$200 = (_$155 ? _$73 : _$45);
    wire [7:0] _$201 = (_$155 ? _$77 : _$12);
    wire _$202 = (_$155 ? _$7 : _$7);
    wire _$203 = (_$198 || _$150);
    wire [7:0] _$204 = (_$198 ? _$199 : _$146);
    wire [7:0] _$205 = (_$198 ? _$200 : _$73);
    wire [7:0] _$206 = (_$198 ? _$201 : _$77);
    wire _$207 = (_$198 ? _$202 : _$28);
    wire _$208 = (_$162 || _$130);
    wire [7:0] _$209 = (_$162 ? _$12 : _$77);
    wire [7:0] _$210 = (_$162 ? _$11 : _$44);
    wire [7:0] _$211 = (_$162 ? _$73 : _$44);
    wire _$212 = (_$162 ? _$28 : _$20);
    wire _$213 = (_$162 ? _$6 : _$28);
    wire _$214 = (_$208 || _$139);
    wire [7:0] _$215 = (_$208 ? _$209 : _$73);
    wire [7:0] _$216 = (_$208 ? _$210 : _$11);
    wire [7:0] _$217 = (_$208 ? _$211 : _$73);
    wire _$218 = (_$208 ? _$212 : _$20);
    wire _$219 = (_$208 ? _$213 : _$6);
    wire _$220 = (_$214 || _$168);
    wire [7:0] _$221 = (_$214 ? _$215 : _$12);
    wire [7:0] _$222 = (_$214 ? _$216 : _$11);
    wire [7:0] _$223 = (_$214 ? _$217 : _$73);
    wire _$224 = (_$214 ? _$218 : _$28);
    wire _$225 = (_$214 ? _$24 : _$28);
    wire _$226 = (_$214 ? _$219 : _$6);
    wire _$227 = (_$156 || _$144);
    wire [7:0] _$228 = (_$156 ? _$146 : _$45);
    wire [7:0] _$229 = (_$156 ? _$73 : _$45);
    wire [7:0] _$230 = (_$156 ? _$77 : _$12);
    wire _$231 = (_$156 ? _$7 : _$7);
    wire _$232 = (_$227 || _$169);
    wire [7:0] _$233 = (_$227 ? _$228 : _$170);
    wire [7:0] _$234 = (_$227 ? _$229 : _$171);
    wire [7:0] _$235 = (_$227 ? _$230 : _$77);
    wire _$236 = (_$227 ? _$231 : _$6);
    reg [2:0] state$;
    always @(posedge clk)
        if (rst) begin
            case (1'b1)
                _$28: state$ <= 3'd0;
            endcase
            reg$wr$5 <= _$28;
            reg$dout$10 <= _$12;
            reg$addr$15 <= _$12;
            reg$rdy$19 <= _$7;
            reg$done$23 <= _$7;
        end else case (state$)
            3'd0: begin
                case (1'b1)
                    _$127: state$ <= 3'd0;
                    _$153: state$ <= 3'd2;
                    _$148: state$ <= 3'd1;
                endcase
                reg$wr$5 <= _$197;
                reg$dout$10 <= _$195;
                reg$addr$15 <= _$194;
                reg$i$43 <= _$196;
            end
            3'd1: begin
                case (1'b1)
                    _$156: state$ <= 3'd2;
                    _$144: state$ <= 3'd3;
                    _$169: state$ <= 3'd1;
                endcase
                reg$wr$5 <= _$236;
                reg$addr$15 <= _$233;
                reg$i$43 <= _$234;
                reg$end$76 <= _$235;
            end
            3'd2: begin
                case (1'b1)
                    _$155: state$ <= 3'd2;
                    _$141: state$ <= 3'd3;
                    _$150: state$ <= 3'd1;
                endcase
                reg$wr$5 <= _$207;
                reg$addr$15 <= _$204;
                reg$i$43 <= _$205;
                reg$end$76 <= _$206;
            end
            3'd3: begin
                case (1'b1)
                    _$28: state$ <= 3'd4;
                endcase
            end
            3'd4: begin
                case (1'b1)
                    _$162: state$ <= 3'd6;
                    _$130: state$ <= 3'd5;
                    _$139: state$ <= 3'd3;
                    _$168: state$ <= 3'd7;
                endcase
                reg$wr$5 <= _$226;
                reg$dout$10 <= _$222;
                reg$addr$15 <= _$221;
                reg$rdy$19 <= _$224;
                reg$done$23 <= _$225;
                reg$i$43 <= _$223;
            end
            3'd5: begin
                case (1'b1)
                    _$160: state$ <= 3'd6;
                    _$138: state$ <= 3'd3;
                    _$166: state$ <= 3'd7;
                endcase
                reg$wr$5 <= _$187;
                reg$addr$15 <= _$182;
                reg$rdy$19 <= _$185;
                reg$done$23 <= _$186;
                reg$i$43 <= _$183;
                reg$end$76 <= _$184;
            end
            3'd6: begin
                case (1'b1)
                    _$158: state$ <= 3'd6;
                    _$164: state$ <= 3'd7;
                endcase
                reg$addr$15 <= _$173;
                reg$done$23 <= _$174;
            end
            3'd7: begin
                case (1'b1)
                    _$28: state$ <= 3'd7;
                endcase
            end
        endcase
endmodule
