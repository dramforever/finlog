module uartrx (clk, rst, in__rx, in__ready, out__data, out__valid);
    input clk;
    input rst;
    input in__rx;
    input in__ready;
    output [7:0] out__data;
    output out__valid;
    reg [7:0] reg__data__6;
    reg reg__valid__11;
    reg [5:0] reg__ctr__22;
    reg [2:0] reg__i__48;
    reg [7:0] reg__cur__52;
    assign out__data = reg__data__6;
    assign out__valid = reg__valid__11;
    wire __0 = in__ready;
    wire __1 = in__rx;
    wire [7:0] __7 = reg__data__6;
    wire [7:0] __8 = 8'd0;
    wire __12 = reg__valid__11;
    wire __13 = 1'b0;
    wire [5:0] __23 = reg__ctr__22;
    wire [5:0] __24 = 6'd0;
    wire [5:0] __35 = 6'd37;
    wire __36 = (__23 != __35);
    wire [5:0] __44 = 6'd1;
    wire [5:0] __45 = (__23 + __44);
    wire [2:0] __49 = reg__i__48;
    wire [2:0] __50 = 3'd0;
    wire [7:0] __53 = reg__cur__52;
    wire [7:0] __54 = 8'd1;
    wire __56 = (__49 != __50);
    wire [7:0] __63 = (__7 | __53);
    wire [7:0] __65 = (__53 + __53);
    wire [2:0] __67 = 3'd1;
    wire [2:0] __68 = (__49 + __67);
    wire [5:0] __71 = 6'd25;
    wire __72 = (__23 != __71);
    wire __84 = 1'b1;
    wire __86 = (! __0);
    wire __100 = (__45 != __35);
    wire __101 = (__84 && __100);
    wire __102 = (! __100);
    wire __103 = (__84 && __102);
    wire __104 = (__45 != __71);
    wire __105 = (__84 && __104);
    wire __106 = (! __104);
    wire __107 = (__84 && __106);
    wire __108 = (__107 && __56);
    wire __109 = (! __56);
    wire __110 = (__107 && __109);
    wire __111 = (__110 && __1);
    wire __112 = (! __1);
    wire __113 = (__110 && __112);
    wire __114 = (__103 && __1);
    wire __115 = (__108 && __1);
    wire __116 = (__103 && __112);
    wire __117 = (__108 && __112);
    wire __118 = (__84 && __86);
    wire __119 = (__111 && __86);
    wire __120 = (! __86);
    wire __121 = (__84 && __120);
    wire __122 = (__111 && __120);
    wire __123 = (__84 && __1);
    wire __124 = (__113 && __1);
    wire __125 = (__84 && __112);
    wire __126 = (__113 && __112);
    wire [7:0] __127 = (__8 | __54);
    wire __128 = (__114 || __116);
    wire [7:0] __129 = (__114 ? __54 : __54);
    wire [5:0] __130 = (__114 ? __45 : __45);
    wire [7:0] __131 = (__114 ? __127 : __8);
    wire [2:0] __132 = (__114 ? __50 : __50);
    wire __133 = (__115 || __117);
    wire [5:0] __134 = (__115 ? __45 : __45);
    wire [7:0] __135 = (__115 ? __63 : __7);
    wire [7:0] __136 = (__129 + __129);
    wire [2:0] __137 = (__132 + __67);
    wire __138 = (__133 || __105);
    wire [7:0] __139 = (__133 ? __65 : __53);
    wire [5:0] __140 = (__133 ? __24 : __45);
    wire [7:0] __141 = (__133 ? __135 : __7);
    wire [2:0] __142 = (__133 ? __68 : __49);
    wire __143 = (__125 || __123);
    wire [5:0] __144 = (__125 ? __24 : __24);
    wire __145 = (__101 || __128);
    wire [7:0] __146 = (__101 ? __53 : __136);
    wire [5:0] __147 = (__101 ? __45 : __24);
    wire [7:0] __148 = (__101 ? __7 : __131);
    wire [2:0] __149 = (__101 ? __49 : __137);
    wire __150 = (__118 || __121);
    wire __151 = (__126 || __119);
    wire __152 = (__126 ? __12 : __84);
    wire [5:0] __153 = (__126 ? __24 : __45);
    wire __154 = (__151 || __138);
    wire __155 = (__151 ? __152 : __12);
    wire [7:0] __156 = (__151 ? __53 : __139);
    wire [5:0] __157 = (__151 ? __153 : __140);
    wire [7:0] __158 = (__151 ? __7 : __141);
    wire [2:0] __159 = (__151 ? __49 : __142);
    wire __160 = (__154 || __124);
    wire __161 = (__154 ? __155 : __12);
    wire [7:0] __162 = (__154 ? __156 : __53);
    wire [5:0] __163 = (__154 ? __157 : __24);
    wire [7:0] __164 = (__154 ? __158 : __7);
    wire [2:0] __165 = (__154 ? __159 : __49);
    wire __166 = (__160 || __122);
    wire __167 = (__160 ? __161 : __84);
    wire [7:0] __168 = (__160 ? __162 : __53);
    wire [5:0] __169 = (__160 ? __163 : __45);
    wire [7:0] __170 = (__160 ? __164 : __7);
    wire [2:0] __171 = (__160 ? __165 : __49);
    wire [5:0] __172 = (__125 ? __24 : __23);
    wire __173 = (__125 ? __13 : __13);
    reg [2:0] state__;
    always @(posedge clk)
        if (rst) begin
            case (1'b1)
                __84: state__ <= 3'd0;
            endcase
            reg__data__6 <= __8;
            reg__valid__11 <= __13;
        end else case (state__)
            3'd0: begin
                case (1'b1)
                    __125: state__ <= 3'd2;
                    __123: state__ <= 3'd1;
                endcase
                reg__ctr__22 <= __144;
            end
            3'd1: begin
                case (1'b1)
                    __125: state__ <= 3'd2;
                    __123: state__ <= 3'd1;
                endcase
                reg__ctr__22 <= __172;
            end
            3'd2: begin
                case (1'b1)
                    __101: state__ <= 3'd2;
                    __128: state__ <= 3'd3;
                endcase
                reg__data__6 <= __148;
                reg__ctr__22 <= __147;
                reg__i__48 <= __149;
                reg__cur__52 <= __146;
            end
            3'd3: begin
                case (1'b1)
                    __126: state__ <= 3'd2;
                    __119: state__ <= 3'd4;
                    __138: state__ <= 3'd3;
                    __124: state__ <= 3'd1;
                    __122: state__ <= 3'd5;
                endcase
                reg__data__6 <= __170;
                reg__valid__11 <= __167;
                reg__ctr__22 <= __169;
                reg__i__48 <= __171;
                reg__cur__52 <= __168;
            end
            3'd4: begin
                case (1'b1)
                    __118: state__ <= 3'd4;
                    __121: state__ <= 3'd5;
                endcase
            end
            3'd5: begin
                case (1'b1)
                    __125: state__ <= 3'd2;
                    __123: state__ <= 3'd1;
                endcase
                reg__valid__11 <= __173;
                reg__ctr__22 <= __144;
            end
        endcase
endmodule
