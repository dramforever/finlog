module lcd (clk, rst, in__data, in__valid, out__rs, out__lcd_out, out__rw, out__ready, out__en);
    input clk;
    input rst;
    input [7:0] in__data;
    input in__valid;
    output out__rs;
    output [7:0] out__lcd_out;
    output out__rw;
    output out__ready;
    output out__en;
    reg reg__ready__6;
    reg reg__en__11;
    reg reg__rs__15;
    reg reg__rw__19;
    reg [7:0] reg__lcd_out__23;
    reg [15:0] reg__ctr__34;
    reg [15:0] reg__ctr__53;
    reg [15:0] reg__ctr__68;
    reg [17:0] reg__ctr__82;
    reg [15:0] reg__ctr__103;
    reg [15:0] reg__ctr__118;
    reg [15:0] reg__ctr__133;
    reg [17:0] reg__ctr__147;
    reg [15:0] reg__ctr__165;
    reg [15:0] reg__ctr__180;
    reg [15:0] reg__ctr__195;
    reg [17:0] reg__ctr__209;
    reg [15:0] reg__ctr__227;
    reg [15:0] reg__ctr__242;
    reg [15:0] reg__ctr__257;
    reg [15:0] reg__ctr__276;
    reg [15:0] reg__ctr__291;
    reg [15:0] reg__ctr__306;
    reg [15:0] reg__ctr__325;
    reg [15:0] reg__ctr__340;
    reg [15:0] reg__ctr__355;
    reg [15:0] reg__ctr__374;
    reg [15:0] reg__ctr__389;
    reg [15:0] reg__ctr__404;
    reg [4:0] reg__count__417;
    reg [7:0] reg__latched__433;
    reg [15:0] reg__ctr__446;
    reg [15:0] reg__ctr__461;
    reg [15:0] reg__ctr__476;
    assign out__rs = reg__rs__15;
    assign out__lcd_out = reg__lcd_out__23;
    assign out__rw = reg__rw__19;
    assign out__ready = reg__ready__6;
    assign out__en = reg__en__11;
    wire [7:0] __0 = in__data;
    wire __1 = in__valid;
    wire __7 = reg__ready__6;
    wire __8 = 1'b0;
    wire __12 = reg__en__11;
    wire __16 = reg__rs__15;
    wire __20 = reg__rw__19;
    wire [7:0] __24 = reg__lcd_out__23;
    wire [7:0] __25 = 8'd0;
    wire [7:0] __31 = 8'd56;
    wire [15:0] __35 = reg__ctr__34;
    wire [15:0] __36 = 16'd0;
    wire [15:0] __38 = 16'd50000;
    wire __39 = (__35 != __38);
    wire [15:0] __47 = 16'd1;
    wire [15:0] __48 = (__35 + __47);
    wire __50 = 1'b1;
    wire [15:0] __54 = reg__ctr__53;
    wire __56 = (__54 != __38);
    wire [15:0] __64 = (__54 + __47);
    wire [15:0] __69 = reg__ctr__68;
    wire __71 = (__69 != __38);
    wire [15:0] __79 = (__69 + __47);
    wire [17:0] __83 = reg__ctr__82;
    wire [17:0] __84 = 18'd0;
    wire [17:0] __86 = 18'd205000;
    wire __87 = (__83 != __86);
    wire [17:0] __95 = 18'd1;
    wire [17:0] __96 = (__83 + __95);
    wire [15:0] __104 = reg__ctr__103;
    wire __106 = (__104 != __38);
    wire [15:0] __114 = (__104 + __47);
    wire [15:0] __119 = reg__ctr__118;
    wire __121 = (__119 != __38);
    wire [15:0] __129 = (__119 + __47);
    wire [15:0] __134 = reg__ctr__133;
    wire __136 = (__134 != __38);
    wire [15:0] __144 = (__134 + __47);
    wire [17:0] __148 = reg__ctr__147;
    wire __150 = (__148 != __86);
    wire [17:0] __158 = (__148 + __95);
    wire [15:0] __166 = reg__ctr__165;
    wire __168 = (__166 != __38);
    wire [15:0] __176 = (__166 + __47);
    wire [15:0] __181 = reg__ctr__180;
    wire __183 = (__181 != __38);
    wire [15:0] __191 = (__181 + __47);
    wire [15:0] __196 = reg__ctr__195;
    wire __198 = (__196 != __38);
    wire [15:0] __206 = (__196 + __47);
    wire [17:0] __210 = reg__ctr__209;
    wire __212 = (__210 != __86);
    wire [17:0] __220 = (__210 + __95);
    wire [15:0] __228 = reg__ctr__227;
    wire __230 = (__228 != __38);
    wire [15:0] __238 = (__228 + __47);
    wire [15:0] __243 = reg__ctr__242;
    wire __245 = (__243 != __38);
    wire [15:0] __253 = (__243 + __47);
    wire [15:0] __258 = reg__ctr__257;
    wire __260 = (__258 != __38);
    wire [15:0] __268 = (__258 + __47);
    wire [7:0] __273 = 8'd1;
    wire [15:0] __277 = reg__ctr__276;
    wire __279 = (__277 != __38);
    wire [15:0] __287 = (__277 + __47);
    wire [15:0] __292 = reg__ctr__291;
    wire __294 = (__292 != __38);
    wire [15:0] __302 = (__292 + __47);
    wire [15:0] __307 = reg__ctr__306;
    wire __309 = (__307 != __38);
    wire [15:0] __317 = (__307 + __47);
    wire [7:0] __322 = 8'd14;
    wire [15:0] __326 = reg__ctr__325;
    wire __328 = (__326 != __38);
    wire [15:0] __336 = (__326 + __47);
    wire [15:0] __341 = reg__ctr__340;
    wire __343 = (__341 != __38);
    wire [15:0] __351 = (__341 + __47);
    wire [15:0] __356 = reg__ctr__355;
    wire __358 = (__356 != __38);
    wire [15:0] __366 = (__356 + __47);
    wire [7:0] __371 = 8'd6;
    wire [15:0] __375 = reg__ctr__374;
    wire __377 = (__375 != __38);
    wire [15:0] __385 = (__375 + __47);
    wire [15:0] __390 = reg__ctr__389;
    wire __392 = (__390 != __38);
    wire [15:0] __400 = (__390 + __47);
    wire [15:0] __405 = reg__ctr__404;
    wire __407 = (__405 != __38);
    wire [15:0] __415 = (__405 + __47);
    wire [4:0] __418 = reg__count__417;
    wire [4:0] __419 = 5'd0;
    wire __424 = (! __1);
    wire [7:0] __434 = reg__latched__433;
    wire [15:0] __447 = reg__ctr__446;
    wire __449 = (__447 != __38);
    wire [15:0] __457 = (__447 + __47);
    wire [15:0] __462 = reg__ctr__461;
    wire __464 = (__462 != __38);
    wire [15:0] __472 = (__462 + __47);
    wire [15:0] __477 = reg__ctr__476;
    wire __479 = (__477 != __38);
    wire [15:0] __487 = (__477 + __47);
    wire __489 = (__114 != __38);
    wire __490 = (__50 && __489);
    wire __491 = (! __489);
    wire __492 = (__50 && __491);
    wire __493 = (__487 != __38);
    wire __494 = (__50 && __493);
    wire __495 = (! __493);
    wire __496 = (__50 && __495);
    wire __497 = (__457 != __38);
    wire __498 = (__50 && __497);
    wire __499 = (! __497);
    wire __500 = (__50 && __499);
    wire __501 = (__472 != __38);
    wire __502 = (__50 && __501);
    wire __503 = (! __501);
    wire __504 = (__50 && __503);
    wire __505 = (__253 != __38);
    wire __506 = (__50 && __505);
    wire __507 = (! __505);
    wire __508 = (__50 && __507);
    wire __509 = (__317 != __38);
    wire __510 = (__50 && __509);
    wire __511 = (! __509);
    wire __512 = (__50 && __511);
    wire __513 = (__220 != __86);
    wire __514 = (__50 && __513);
    wire __515 = (! __513);
    wire __516 = (__50 && __515);
    wire __517 = (__268 != __38);
    wire __518 = (__50 && __517);
    wire __519 = (! __517);
    wire __520 = (__50 && __519);
    wire __521 = (__415 != __38);
    wire __522 = (__50 && __521);
    wire __523 = (! __521);
    wire __524 = (__50 && __523);
    wire __525 = (__191 != __38);
    wire __526 = (__50 && __525);
    wire __527 = (! __525);
    wire __528 = (__50 && __527);
    wire __529 = (__287 != __38);
    wire __530 = (__50 && __529);
    wire __531 = (! __529);
    wire __532 = (__50 && __531);
    wire __533 = (__48 != __38);
    wire __534 = (__50 && __533);
    wire __535 = (! __533);
    wire __536 = (__50 && __535);
    wire __537 = (__96 != __86);
    wire __538 = (__50 && __537);
    wire __539 = (! __537);
    wire __540 = (__50 && __539);
    wire __541 = (__351 != __38);
    wire __542 = (__50 && __541);
    wire __543 = (! __541);
    wire __544 = (__50 && __543);
    wire __545 = (__79 != __38);
    wire __546 = (__50 && __545);
    wire __547 = (! __545);
    wire __548 = (__50 && __547);
    wire __549 = (__158 != __86);
    wire __550 = (__50 && __549);
    wire __551 = (! __549);
    wire __552 = (__50 && __551);
    wire __553 = (__206 != __38);
    wire __554 = (__50 && __553);
    wire __555 = (! __553);
    wire __556 = (__50 && __555);
    wire __557 = (__238 != __38);
    wire __558 = (__50 && __557);
    wire __559 = (! __557);
    wire __560 = (__50 && __559);
    wire __561 = (__302 != __38);
    wire __562 = (__50 && __561);
    wire __563 = (! __561);
    wire __564 = (__50 && __563);
    wire __565 = (__366 != __38);
    wire __566 = (__50 && __565);
    wire __567 = (! __565);
    wire __568 = (__50 && __567);
    wire __569 = (__129 != __38);
    wire __570 = (__50 && __569);
    wire __571 = (! __569);
    wire __572 = (__50 && __571);
    wire __573 = (__385 != __38);
    wire __574 = (__50 && __573);
    wire __575 = (! __573);
    wire __576 = (__50 && __575);
    wire __577 = (__144 != __38);
    wire __578 = (__50 && __577);
    wire __579 = (! __577);
    wire __580 = (__50 && __579);
    wire __581 = (__400 != __38);
    wire __582 = (__50 && __581);
    wire __583 = (! __581);
    wire __584 = (__50 && __583);
    wire __585 = (__176 != __38);
    wire __586 = (__50 && __585);
    wire __587 = (! __585);
    wire __588 = (__50 && __587);
    wire __589 = (__64 != __38);
    wire __590 = (__50 && __589);
    wire __591 = (! __589);
    wire __592 = (__50 && __591);
    wire __593 = (__336 != __38);
    wire __594 = (__50 && __593);
    wire __595 = (! __593);
    wire __596 = (__50 && __595);
    wire __597 = (__496 && __424);
    wire __598 = (__524 && __424);
    wire __599 = (__50 && __424);
    wire __600 = (! __424);
    wire __601 = (__496 && __600);
    wire __602 = (__524 && __600);
    wire __603 = (__50 && __600);
    wire __604 = (__494 || __601);
    wire __605 = (__494 ? __7 : __50);
    wire [15:0] __606 = (__494 ? __487 : __487);
    wire [7:0] __607 = (__494 ? __434 : __0);
    wire __608 = (__604 || __597);
    wire __609 = (__604 ? __605 : __50);
    wire [15:0] __610 = (__604 ? __606 : __487);
    wire [7:0] __611 = (__604 ? __607 : __434);
    wire __612 = (__504 || __502);
    wire [15:0] __613 = (__504 ? __472 : __472);
    wire __614 = (__504 ? __8 : __12);
    wire [15:0] __615 = (__504 ? __36 : __477);
    wire __616 = (__500 || __498);
    wire [15:0] __617 = (__500 ? __36 : __462);
    wire __618 = (__500 ? __50 : __12);
    wire [15:0] __619 = (__500 ? __457 : __457);
    wire __620 = (__518 || __520);
    wire [15:0] __621 = (__518 ? __268 : __268);
    wire __622 = (__518 ? __20 : __8);
    wire [15:0] __623 = (__518 ? __277 : __36);
    wire [7:0] __624 = (__518 ? __24 : __273);
    wire __625 = (__518 ? __16 : __8);
    wire __626 = (__514 || __516);
    wire [17:0] __627 = (__514 ? __220 : __220);
    wire [15:0] __628 = (__514 ? __228 : __36);
    wire __629 = (__514 ? __20 : __8);
    wire [7:0] __630 = (__514 ? __24 : __31);
    wire __631 = (__514 ? __16 : __8);
    wire __632 = (__510 || __512);
    wire __633 = (__510 ? __20 : __8);
    wire [15:0] __634 = (__510 ? __317 : __317);
    wire [15:0] __635 = (__510 ? __326 : __36);
    wire [7:0] __636 = (__510 ? __24 : __322);
    wire __637 = (__510 ? __16 : __8);
    wire __638 = (__508 || __506);
    wire [15:0] __639 = (__508 ? __36 : __258);
    wire [15:0] __640 = (__508 ? __253 : __253);
    wire __641 = (__508 ? __8 : __12);
    wire __642 = (__564 || __562);
    wire [15:0] __643 = (__564 ? __302 : __302);
    wire [15:0] __644 = (__564 ? __36 : __307);
    wire __645 = (__564 ? __8 : __12);
    wire __646 = (__566 || __568);
    wire __647 = (__566 ? __20 : __8);
    wire [15:0] __648 = (__566 ? __366 : __366);
    wire [15:0] __649 = (__566 ? __375 : __36);
    wire [7:0] __650 = (__566 ? __24 : __371);
    wire __651 = (__566 ? __16 : __8);
    wire __652 = (__550 || __552);
    wire __653 = (__550 ? __20 : __8);
    wire [17:0] __654 = (__550 ? __158 : __158);
    wire [15:0] __655 = (__550 ? __166 : __36);
    wire [7:0] __656 = (__550 ? __24 : __31);
    wire __657 = (__550 ? __16 : __8);
    wire __658 = (__556 || __554);
    wire [17:0] __659 = (__556 ? __84 : __210);
    wire [15:0] __660 = (__556 ? __206 : __206);
    wire __661 = (__560 || __558);
    wire [15:0] __662 = (__560 ? __238 : __238);
    wire [15:0] __663 = (__560 ? __36 : __243);
    wire __664 = (__560 ? __50 : __12);
    wire __665 = (__532 || __530);
    wire [15:0] __666 = (__532 ? __36 : __292);
    wire [15:0] __667 = (__532 ? __287 : __287);
    wire __668 = (__532 ? __50 : __12);
    wire __669 = (__534 || __536);
    wire [15:0] __670 = (__534 ? __48 : __48);
    wire [15:0] __671 = (__534 ? __54 : __36);
    wire __672 = (__534 ? __12 : __50);
    wire __673 = (__546 || __548);
    wire [17:0] __674 = (__546 ? __83 : __84);
    wire [15:0] __675 = (__546 ? __79 : __79);
    wire __676 = (__538 || __540);
    wire __677 = (__538 ? __20 : __8);
    wire [17:0] __678 = (__538 ? __96 : __96);
    wire [15:0] __679 = (__538 ? __104 : __36);
    wire [7:0] __680 = (__538 ? __24 : __31);
    wire __681 = (__538 ? __16 : __8);
    wire __682 = (__544 || __542);
    wire [15:0] __683 = (__544 ? __36 : __356);
    wire [15:0] __684 = (__544 ? __351 : __351);
    wire __685 = (__544 ? __8 : __12);
    wire __686 = (__602 || __522);
    wire __687 = (__602 ? __50 : __7);
    wire [15:0] __688 = (__602 ? __415 : __415);
    wire [7:0] __689 = (__602 ? __0 : __434);
    wire [4:0] __690 = (__602 ? __419 : __418);
    wire __691 = (__686 || __598);
    wire __692 = (__686 ? __687 : __50);
    wire [15:0] __693 = (__686 ? __688 : __415);
    wire [7:0] __694 = (__686 ? __689 : __434);
    wire [4:0] __695 = (__686 ? __690 : __419);
    wire __696 = (__528 || __526);
    wire [15:0] __697 = (__528 ? __36 : __196);
    wire [15:0] __698 = (__528 ? __191 : __191);
    wire __699 = (__528 ? __8 : __12);
    wire __700 = (__592 || __590);
    wire [15:0] __701 = (__592 ? __64 : __64);
    wire [15:0] __702 = (__592 ? __36 : __69);
    wire __703 = (__592 ? __8 : __12);
    wire __704 = (__596 || __594);
    wire [15:0] __705 = (__596 ? __336 : __336);
    wire [15:0] __706 = (__596 ? __36 : __341);
    wire __707 = (__596 ? __50 : __12);
    wire __708 = (__580 || __578);
    wire [17:0] __709 = (__580 ? __84 : __148);
    wire [15:0] __710 = (__580 ? __144 : __144);
    wire __711 = (__584 || __582);
    wire [15:0] __712 = (__584 ? __400 : __400);
    wire [15:0] __713 = (__584 ? __36 : __405);
    wire __714 = (__584 ? __8 : __12);
    wire __715 = (__588 || __586);
    wire [15:0] __716 = (__588 ? __176 : __176);
    wire [15:0] __717 = (__588 ? __36 : __181);
    wire __718 = (__588 ? __50 : __12);
    wire __719 = (__603 || __599);
    wire [7:0] __720 = (__603 ? __0 : __434);
    wire __721 = (__572 || __570);
    wire [15:0] __722 = (__572 ? __36 : __134);
    wire [15:0] __723 = (__572 ? __129 : __129);
    wire __724 = (__572 ? __8 : __12);
    wire __725 = (__576 || __574);
    wire [15:0] __726 = (__576 ? __36 : __390);
    wire [15:0] __727 = (__576 ? __385 : __385);
    wire __728 = (__576 ? __50 : __12);
    wire __729 = (__492 || __490);
    wire [15:0] __730 = (__492 ? __114 : __114);
    wire [15:0] __731 = (__492 ? __36 : __119);
    wire __732 = (__492 ? __50 : __12);
    reg [4:0] state__;
    always @(posedge clk)
        if (rst) begin
            case (1'b1)
                __50: state__ <= 5'd0;
            endcase
            reg__ready__6 <= __8;
            reg__en__11 <= __8;
            reg__rs__15 <= __8;
            reg__rw__19 <= __8;
            reg__lcd_out__23 <= __31;
            reg__ctr__34 <= __36;
        end else case (state__)
            5'd0: begin
                case (1'b1)
                    __534: state__ <= 5'd0;
                    __536: state__ <= 5'd1;
                endcase
                reg__en__11 <= __672;
                reg__ctr__34 <= __670;
                reg__ctr__53 <= __671;
            end
            5'd1: begin
                case (1'b1)
                    __592: state__ <= 5'd2;
                    __590: state__ <= 5'd1;
                endcase
                reg__en__11 <= __703;
                reg__ctr__53 <= __701;
                reg__ctr__68 <= __702;
            end
            5'd2: begin
                case (1'b1)
                    __546: state__ <= 5'd2;
                    __548: state__ <= 5'd3;
                endcase
                reg__ctr__68 <= __675;
                reg__ctr__82 <= __674;
            end
            5'd3: begin
                case (1'b1)
                    __538: state__ <= 5'd3;
                    __540: state__ <= 5'd4;
                endcase
                reg__rs__15 <= __681;
                reg__rw__19 <= __677;
                reg__lcd_out__23 <= __680;
                reg__ctr__82 <= __678;
                reg__ctr__103 <= __679;
            end
            5'd4: begin
                case (1'b1)
                    __492: state__ <= 5'd5;
                    __490: state__ <= 5'd4;
                endcase
                reg__en__11 <= __732;
                reg__ctr__103 <= __730;
                reg__ctr__118 <= __731;
            end
            5'd5: begin
                case (1'b1)
                    __572: state__ <= 5'd6;
                    __570: state__ <= 5'd5;
                endcase
                reg__en__11 <= __724;
                reg__ctr__118 <= __723;
                reg__ctr__133 <= __722;
            end
            5'd6: begin
                case (1'b1)
                    __580: state__ <= 5'd7;
                    __578: state__ <= 5'd6;
                endcase
                reg__ctr__133 <= __710;
                reg__ctr__147 <= __709;
            end
            5'd7: begin
                case (1'b1)
                    __550: state__ <= 5'd7;
                    __552: state__ <= 5'd8;
                endcase
                reg__rs__15 <= __657;
                reg__rw__19 <= __653;
                reg__lcd_out__23 <= __656;
                reg__ctr__147 <= __654;
                reg__ctr__165 <= __655;
            end
            5'd8: begin
                case (1'b1)
                    __588: state__ <= 5'd9;
                    __586: state__ <= 5'd8;
                endcase
                reg__en__11 <= __718;
                reg__ctr__165 <= __716;
                reg__ctr__180 <= __717;
            end
            5'd9: begin
                case (1'b1)
                    __528: state__ <= 5'd10;
                    __526: state__ <= 5'd9;
                endcase
                reg__en__11 <= __699;
                reg__ctr__180 <= __698;
                reg__ctr__195 <= __697;
            end
            5'd10: begin
                case (1'b1)
                    __556: state__ <= 5'd11;
                    __554: state__ <= 5'd10;
                endcase
                reg__ctr__195 <= __660;
                reg__ctr__209 <= __659;
            end
            5'd11: begin
                case (1'b1)
                    __514: state__ <= 5'd11;
                    __516: state__ <= 5'd12;
                endcase
                reg__rs__15 <= __631;
                reg__rw__19 <= __629;
                reg__lcd_out__23 <= __630;
                reg__ctr__209 <= __627;
                reg__ctr__227 <= __628;
            end
            5'd12: begin
                case (1'b1)
                    __560: state__ <= 5'd13;
                    __558: state__ <= 5'd12;
                endcase
                reg__en__11 <= __664;
                reg__ctr__227 <= __662;
                reg__ctr__242 <= __663;
            end
            5'd13: begin
                case (1'b1)
                    __508: state__ <= 5'd14;
                    __506: state__ <= 5'd13;
                endcase
                reg__en__11 <= __641;
                reg__ctr__242 <= __640;
                reg__ctr__257 <= __639;
            end
            5'd14: begin
                case (1'b1)
                    __518: state__ <= 5'd14;
                    __520: state__ <= 5'd15;
                endcase
                reg__rs__15 <= __625;
                reg__rw__19 <= __622;
                reg__lcd_out__23 <= __624;
                reg__ctr__257 <= __621;
                reg__ctr__276 <= __623;
            end
            5'd15: begin
                case (1'b1)
                    __532: state__ <= 5'd16;
                    __530: state__ <= 5'd15;
                endcase
                reg__en__11 <= __668;
                reg__ctr__276 <= __667;
                reg__ctr__291 <= __666;
            end
            5'd16: begin
                case (1'b1)
                    __564: state__ <= 5'd17;
                    __562: state__ <= 5'd16;
                endcase
                reg__en__11 <= __645;
                reg__ctr__291 <= __643;
                reg__ctr__306 <= __644;
            end
            5'd17: begin
                case (1'b1)
                    __510: state__ <= 5'd17;
                    __512: state__ <= 5'd18;
                endcase
                reg__rs__15 <= __637;
                reg__rw__19 <= __633;
                reg__lcd_out__23 <= __636;
                reg__ctr__306 <= __634;
                reg__ctr__325 <= __635;
            end
            5'd18: begin
                case (1'b1)
                    __596: state__ <= 5'd19;
                    __594: state__ <= 5'd18;
                endcase
                reg__en__11 <= __707;
                reg__ctr__325 <= __705;
                reg__ctr__340 <= __706;
            end
            5'd19: begin
                case (1'b1)
                    __544: state__ <= 5'd20;
                    __542: state__ <= 5'd19;
                endcase
                reg__en__11 <= __685;
                reg__ctr__340 <= __684;
                reg__ctr__355 <= __683;
            end
            5'd20: begin
                case (1'b1)
                    __566: state__ <= 5'd20;
                    __568: state__ <= 5'd21;
                endcase
                reg__rs__15 <= __651;
                reg__rw__19 <= __647;
                reg__lcd_out__23 <= __650;
                reg__ctr__355 <= __648;
                reg__ctr__374 <= __649;
            end
            5'd21: begin
                case (1'b1)
                    __576: state__ <= 5'd22;
                    __574: state__ <= 5'd21;
                endcase
                reg__en__11 <= __728;
                reg__ctr__374 <= __727;
                reg__ctr__389 <= __726;
            end
            5'd22: begin
                case (1'b1)
                    __584: state__ <= 5'd23;
                    __582: state__ <= 5'd22;
                endcase
                reg__en__11 <= __714;
                reg__ctr__389 <= __712;
                reg__ctr__404 <= __713;
            end
            5'd23: begin
                case (1'b1)
                    __602: state__ <= 5'd25;
                    __522: state__ <= 5'd23;
                    __598: state__ <= 5'd24;
                endcase
                reg__ready__6 <= __692;
                reg__ctr__404 <= __693;
                reg__count__417 <= __695;
                reg__latched__433 <= __694;
            end
            5'd24: begin
                case (1'b1)
                    __603: state__ <= 5'd25;
                    __599: state__ <= 5'd24;
                endcase
                reg__latched__433 <= __720;
            end
            5'd25: begin
                case (1'b1)
                    __50: state__ <= 5'd26;
                endcase
                reg__ready__6 <= __8;
                reg__rs__15 <= __50;
                reg__rw__19 <= __8;
                reg__lcd_out__23 <= __434;
                reg__ctr__446 <= __36;
            end
            5'd26: begin
                case (1'b1)
                    __500: state__ <= 5'd27;
                    __498: state__ <= 5'd26;
                endcase
                reg__en__11 <= __618;
                reg__ctr__446 <= __619;
                reg__ctr__461 <= __617;
            end
            5'd27: begin
                case (1'b1)
                    __504: state__ <= 5'd28;
                    __502: state__ <= 5'd27;
                endcase
                reg__en__11 <= __614;
                reg__ctr__461 <= __613;
                reg__ctr__476 <= __615;
            end
            5'd28: begin
                case (1'b1)
                    __494: state__ <= 5'd28;
                    __601: state__ <= 5'd25;
                    __597: state__ <= 5'd24;
                endcase
                reg__ready__6 <= __609;
                reg__latched__433 <= __611;
                reg__ctr__476 <= __610;
            end
        endcase
endmodule
