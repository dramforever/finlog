module sieve (clk, rst, in__din, out__wr, out__done, out__addr, out__rdy, out__dout);
    input clk;
    input rst;
    input [7:0] in__din;
    output out__wr;
    output out__done;
    output [7:0] out__addr;
    output out__rdy;
    output [7:0] out__dout;
    reg reg__wr__5;
    reg [7:0] reg__dout__10;
    reg [7:0] reg__addr__15;
    reg reg__rdy__19;
    reg reg__done__23;
    reg [7:0] reg__i__43;
    reg [7:0] reg__end__76;
    assign out__wr = reg__wr__5;
    assign out__done = reg__done__23;
    assign out__addr = reg__addr__15;
    assign out__rdy = reg__rdy__19;
    assign out__dout = reg__dout__10;
    wire [7:0] __0 = in__din;
    wire __6 = reg__wr__5;
    wire __7 = 1'b0;
    wire [7:0] __11 = reg__dout__10;
    wire [7:0] __12 = 8'd0;
    wire [7:0] __16 = reg__addr__15;
    wire __20 = reg__rdy__19;
    wire __24 = reg__done__23;
    wire __28 = 1'b1;
    wire [7:0] __31 = 8'd100;
    wire __32 = (__16 <= __31);
    wire [7:0] __40 = 8'd1;
    wire [7:0] __41 = (__16 + __40);
    wire [7:0] __44 = reg__i__43;
    wire [7:0] __45 = 8'd2;
    wire __48 = (__44 <= __31);
    wire [7:0] __52 = (__44 + __44);
    wire [7:0] __64 = (__16 + __44);
    wire [7:0] __73 = (__44 + __40);
    wire [7:0] __77 = reg__end__76;
    wire __94 = (! __0);
    wire [7:0] __104 = (__77 + __40);
    wire __109 = (__16 < __77);
    wire __126 = (__41 <= __31);
    wire __127 = (__28 && __126);
    wire __128 = (! __126);
    wire __129 = (__28 && __128);
    wire __130 = (__28 && __94);
    wire __131 = (! __94);
    wire __132 = (__28 && __131);
    wire __133 = (__64 <= __31);
    wire __134 = (__28 && __133);
    wire __135 = (! __133);
    wire __136 = (__28 && __135);
    wire __137 = (__73 <= __31);
    wire __138 = (__28 && __137);
    wire __139 = (__132 && __137);
    wire __140 = (! __137);
    wire __141 = (__28 && __140);
    wire __142 = (__132 && __140);
    wire __143 = (__136 && __137);
    wire __144 = (__136 && __140);
    wire [7:0] __145 = (__45 + __45);
    wire [7:0] __146 = (__73 + __73);
    wire __147 = (__145 <= __31);
    wire __148 = (__129 && __147);
    wire __149 = (__146 <= __31);
    wire __150 = (__138 && __149);
    wire __151 = (__143 && __149);
    wire __152 = (! __147);
    wire __153 = (__129 && __152);
    wire __154 = (! __149);
    wire __155 = (__138 && __154);
    wire __156 = (__143 && __154);
    wire __157 = (__41 < __77);
    wire __158 = (__28 && __157);
    wire __159 = (__12 < __104);
    wire __160 = (__141 && __159);
    wire __161 = (__12 < __77);
    wire __162 = (__142 && __161);
    wire __163 = (! __157);
    wire __164 = (__28 && __163);
    wire __165 = (! __159);
    wire __166 = (__141 && __165);
    wire __167 = (! __161);
    wire __168 = (__142 && __167);
    wire __169 = (__151 || __134);
    wire [7:0] __170 = (__151 ? __146 : __64);
    wire [7:0] __171 = (__151 ? __73 : __44);
    wire __172 = (__158 || __164);
    wire [7:0] __173 = (__158 ? __41 : __41);
    wire __174 = (__158 ? __24 : __28);
    wire __175 = (__160 || __138);
    wire [7:0] __176 = (__160 ? __12 : __73);
    wire [7:0] __177 = (__160 ? __73 : __73);
    wire [7:0] __178 = (__160 ? __104 : __104);
    wire __179 = (__160 ? __28 : __20);
    wire __180 = (__160 ? __7 : __7);
    wire __181 = (__175 || __166);
    wire [7:0] __182 = (__175 ? __176 : __12);
    wire [7:0] __183 = (__175 ? __177 : __73);
    wire [7:0] __184 = (__175 ? __178 : __104);
    wire __185 = (__175 ? __179 : __28);
    wire __186 = (__175 ? __24 : __28);
    wire __187 = (__175 ? __180 : __7);
    wire __188 = (__127 || __153);
    wire [7:0] __189 = (__127 ? __41 : __145);
    wire [7:0] __190 = (__127 ? __11 : __40);
    wire [7:0] __191 = (__127 ? __44 : __45);
    wire __192 = (__127 ? __6 : __7);
    wire __193 = (__188 || __148);
    wire [7:0] __194 = (__188 ? __189 : __145);
    wire [7:0] __195 = (__188 ? __190 : __40);
    wire [7:0] __196 = (__188 ? __191 : __45);
    wire __197 = (__188 ? __192 : __6);
    wire __198 = (__155 || __141);
    wire [7:0] __199 = (__155 ? __146 : __45);
    wire [7:0] __200 = (__155 ? __73 : __45);
    wire [7:0] __201 = (__155 ? __77 : __12);
    wire __202 = (__155 ? __7 : __7);
    wire __203 = (__198 || __150);
    wire [7:0] __204 = (__198 ? __199 : __146);
    wire [7:0] __205 = (__198 ? __200 : __73);
    wire [7:0] __206 = (__198 ? __201 : __77);
    wire __207 = (__198 ? __202 : __28);
    wire __208 = (__162 || __130);
    wire [7:0] __209 = (__162 ? __12 : __77);
    wire [7:0] __210 = (__162 ? __11 : __44);
    wire [7:0] __211 = (__162 ? __73 : __44);
    wire __212 = (__162 ? __28 : __20);
    wire __213 = (__162 ? __6 : __28);
    wire __214 = (__208 || __139);
    wire [7:0] __215 = (__208 ? __209 : __73);
    wire [7:0] __216 = (__208 ? __210 : __11);
    wire [7:0] __217 = (__208 ? __211 : __73);
    wire __218 = (__208 ? __212 : __20);
    wire __219 = (__208 ? __213 : __6);
    wire __220 = (__214 || __168);
    wire [7:0] __221 = (__214 ? __215 : __12);
    wire [7:0] __222 = (__214 ? __216 : __11);
    wire [7:0] __223 = (__214 ? __217 : __73);
    wire __224 = (__214 ? __218 : __28);
    wire __225 = (__214 ? __24 : __28);
    wire __226 = (__214 ? __219 : __6);
    wire __227 = (__156 || __144);
    wire [7:0] __228 = (__156 ? __146 : __45);
    wire [7:0] __229 = (__156 ? __73 : __45);
    wire [7:0] __230 = (__156 ? __77 : __12);
    wire __231 = (__156 ? __7 : __7);
    wire __232 = (__227 || __169);
    wire [7:0] __233 = (__227 ? __228 : __170);
    wire [7:0] __234 = (__227 ? __229 : __171);
    wire [7:0] __235 = (__227 ? __230 : __77);
    wire __236 = (__227 ? __231 : __6);
    reg [2:0] state__;
    always @(posedge clk)
        if (rst) begin
            case (1'b1)
                __28: state__ <= 3'd0;
            endcase
            reg__wr__5 <= __28;
            reg__dout__10 <= __12;
            reg__addr__15 <= __12;
            reg__rdy__19 <= __7;
            reg__done__23 <= __7;
        end else case (state__)
            3'd0: begin
                case (1'b1)
                    __127: state__ <= 3'd0;
                    __153: state__ <= 3'd2;
                    __148: state__ <= 3'd1;
                endcase
                reg__wr__5 <= __197;
                reg__dout__10 <= __195;
                reg__addr__15 <= __194;
                reg__i__43 <= __196;
            end
            3'd1: begin
                case (1'b1)
                    __156: state__ <= 3'd2;
                    __144: state__ <= 3'd3;
                    __169: state__ <= 3'd1;
                endcase
                reg__wr__5 <= __236;
                reg__addr__15 <= __233;
                reg__i__43 <= __234;
                reg__end__76 <= __235;
            end
            3'd2: begin
                case (1'b1)
                    __155: state__ <= 3'd2;
                    __141: state__ <= 3'd3;
                    __150: state__ <= 3'd1;
                endcase
                reg__wr__5 <= __207;
                reg__addr__15 <= __204;
                reg__i__43 <= __205;
                reg__end__76 <= __206;
            end
            3'd3: begin
                case (1'b1)
                    __28: state__ <= 3'd4;
                endcase
            end
            3'd4: begin
                case (1'b1)
                    __162: state__ <= 3'd6;
                    __130: state__ <= 3'd5;
                    __139: state__ <= 3'd3;
                    __168: state__ <= 3'd7;
                endcase
                reg__wr__5 <= __226;
                reg__dout__10 <= __222;
                reg__addr__15 <= __221;
                reg__rdy__19 <= __224;
                reg__done__23 <= __225;
                reg__i__43 <= __223;
            end
            3'd5: begin
                case (1'b1)
                    __160: state__ <= 3'd6;
                    __138: state__ <= 3'd3;
                    __166: state__ <= 3'd7;
                endcase
                reg__wr__5 <= __187;
                reg__addr__15 <= __182;
                reg__rdy__19 <= __185;
                reg__done__23 <= __186;
                reg__i__43 <= __183;
                reg__end__76 <= __184;
            end
            3'd6: begin
                case (1'b1)
                    __158: state__ <= 3'd6;
                    __164: state__ <= 3'd7;
                endcase
                reg__addr__15 <= __173;
                reg__done__23 <= __174;
            end
            3'd7: begin
                case (1'b1)
                    __28: state__ <= 3'd7;
                endcase
            end
        endcase
endmodule
